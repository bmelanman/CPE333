module cache_structure (
    input logic clk,
    input logic rst
);


endmodule : cache_structure
