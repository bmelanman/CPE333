
module top;

    cam_if itf ();
    testbench tb (.*);
    grader gdr (.*);

endmodule : top
